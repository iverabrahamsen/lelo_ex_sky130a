magic
tech sky130A
magscale 1 2
timestamp 1768564347
<< locali >>
rect 193 1960 419 2040
rect -96 -200 96 152
rect 1056 -200 1248 152
rect -200 -207 1400 -200
rect -200 -387 294 -207
rect 474 -387 1400 -207
rect -200 -400 1400 -387
<< viali >>
rect 294 -387 474 -207
<< metal1 >>
rect 160 43 224 3304
rect 288 -207 480 3888
rect 672 3832 864 4007
rect 672 3640 1154 3832
rect 672 3252 864 3640
rect 966 3063 1151 3640
rect 672 2871 1151 3063
rect 672 1175 864 1454
rect 966 1175 1151 2871
rect 672 983 1151 1175
rect 966 386 1151 983
rect 698 201 1151 386
rect 672 40 864 120
rect 288 -387 294 -207
rect 474 -387 480 -207
rect 288 -399 480 -387
use JNWATR_NCH_4C5F0  xo0<0> ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 0
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo0<1>
timestamp 1740610800
transform 1 0 0 0 1 800
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1<0>
timestamp 1740610800
transform 1 0 0 0 1 2400
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1<1>
timestamp 1740610800
transform 1 0 0 0 1 3200
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1
timestamp 1740610800
transform 1 0 0 0 1 1600
box -184 -128 1336 928
<< labels >>
flabel metal1 s 288 600 480 680 0 FreeSans 400 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal1 s 160 360 224 440 0 FreeSans 400 0 0 0 IBPS_5U
port 2 nsew signal bidirectional
flabel metal1 s 672 40 864 120 0 FreeSans 400 0 0 0 IBNS_20U
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 4000
<< end >>
